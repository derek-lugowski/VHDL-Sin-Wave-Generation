library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity volt2dist is 
	port(
		volt		: in	std_logic_vector(11 downto 0);
		dist		: out	std_logic_vector(12 downto 0)
		);
end volt2dist;

architecture lookupTable of volt2dist is


type rom is array (0 to 4095) of integer;

constant table: rom:=(       --distance (cm * 100)
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(3292),
(3281),
(3271),
(3261),
(3250),
(3240),
(3230),
(3220),
(3210),
(3200),
(3190),
(3180),
(3170),
(3160),
(3151),
(3141),
(3132),
(3122),
(3113),
(3103),
(3094),
(3084),
(3075),
(3066),
(3057),
(3048),
(3039),
(3030),
(3021),
(3012),
(3003),
(2994),
(2986),
(2977),
(2968),
(2960),
(2951),
(2943),
(2934),
(2926),
(2917),
(2909),
(2901),
(2893),
(2884),
(2876),
(2868),
(2860),
(2852),
(2844),
(2836),
(2828),
(2821),
(2813),
(2805),
(2797),
(2790),
(2782),
(2775),
(2767),
(2759),
(2752),
(2745),
(2737),
(2730),
(2723),
(2715),
(2708),
(2701),
(2694),
(2687),
(2679),
(2672),
(2665),
(2658),
(2651),
(2645),
(2638),
(2631),
(2624),
(2617),
(2611),
(2604),
(2597),
(2591),
(2584),
(2577),
(2571),
(2564),
(2558),
(2551),
(2545),
(2539),
(2532),
(2526),
(2520),
(2513),
(2507),
(2501),
(2495),
(2489),
(2483),
(2476),
(2470),
(2464),
(2458),
(2452),
(2446),
(2441),
(2435),
(2429),
(2423),
(2417),
(2411),
(2406),
(2400),
(2394),
(2389),
(2383),
(2377),
(2372),
(2366),
(2361),
(2355),
(2350),
(2344),
(2339),
(2333),
(2328),
(2322),
(2317),
(2312),
(2306),
(2301),
(2296),
(2291),
(2285),
(2280),
(2275),
(2270),
(2265),
(2260),
(2255),
(2250),
(2245),
(2240),
(2235),
(2230),
(2225),
(2220),
(2215),
(2210),
(2205),
(2200),
(2195),
(2191),
(2186),
(2181),
(2176),
(2172),
(2167),
(2162),
(2158),
(2153),
(2148),
(2144),
(2139),
(2135),
(2130),
(2126),
(2121),
(2117),
(2112),
(2108),
(2103),
(2099),
(2094),
(2090),
(2086),
(2081),
(2077),
(2073),
(2068),
(2064),
(2060),
(2056),
(2051),
(2047),
(2043),
(2039),
(2035),
(2031),
(2026),
(2022),
(2018),
(2014),
(2010),
(2006),
(2002),
(1998),
(1994),
(1990),
(1986),
(1982),
(1978),
(1974),
(1970),
(1966),
(1963),
(1959),
(1955),
(1951),
(1947),
(1943),
(1940),
(1936),
(1932),
(1928),
(1925),
(1921),
(1917),
(1913),
(1910),
(1906),
(1902),
(1899),
(1895),
(1892),
(1888),
(1884),
(1881),
(1877),
(1874),
(1870),
(1867),
(1863),
(1860),
(1856),
(1853),
(1849),
(1846),
(1842),
(1839),
(1836),
(1832),
(1829),
(1825),
(1822),
(1819),
(1815),
(1812),
(1809),
(1805),
(1802),
(1799),
(1796),
(1792),
(1789),
(1786),
(1783),
(1779),
(1776),
(1773),
(1770),
(1767),
(1764),
(1760),
(1757),
(1754),
(1751),
(1748),
(1745),
(1742),
(1739),
(1736),
(1733),
(1730),
(1727),
(1724),
(1720),
(1717),
(1715),
(1712),
(1709),
(1706),
(1703),
(1700),
(1697),
(1694),
(1691),
(1688),
(1685),
(1682),
(1679),
(1677),
(1674),
(1671),
(1668),
(1665),
(1662),
(1660),
(1657),
(1654),
(1651),
(1649),
(1646),
(1643),
(1640),
(1638),
(1635),
(1632),
(1629),
(1627),
(1624),
(1621),
(1619),
(1616),
(1613),
(1611),
(1608),
(1605),
(1603),
(1600),
(1598),
(1595),
(1592),
(1590),
(1587),
(1585),
(1582),
(1580),
(1577),
(1575),
(1572),
(1569),
(1567),
(1564),
(1562),
(1559),
(1557),
(1555),
(1552),
(1550),
(1547),
(1545),
(1542),
(1540),
(1537),
(1535),
(1533),
(1530),
(1528),
(1525),
(1523),
(1521),
(1518),
(1516),
(1514),
(1511),
(1509),
(1507),
(1504),
(1502),
(1500),
(1497),
(1495),
(1493),
(1491),
(1488),
(1486),
(1484),
(1482),
(1479),
(1477),
(1475),
(1473),
(1470),
(1468),
(1466),
(1464),
(1462),
(1459),
(1457),
(1455),
(1453),
(1451),
(1449),
(1446),
(1444),
(1442),
(1440),
(1438),
(1436),
(1434),
(1432),
(1429),
(1427),
(1425),
(1423),
(1421),
(1419),
(1417),
(1415),
(1413),
(1411),
(1409),
(1407),
(1405),
(1403),
(1401),
(1399),
(1397),
(1395),
(1393),
(1391),
(1389),
(1387),
(1385),
(1383),
(1381),
(1379),
(1377),
(1375),
(1373),
(1371),
(1369),
(1367),
(1365),
(1363),
(1361),
(1360),
(1358),
(1356),
(1354),
(1352),
(1350),
(1348),
(1346),
(1344),
(1343),
(1341),
(1339),
(1337),
(1335),
(1333),
(1332),
(1330),
(1328),
(1326),
(1324),
(1322),
(1321),
(1319),
(1317),
(1315),
(1313),
(1312),
(1310),
(1308),
(1306),
(1305),
(1303),
(1301),
(1299),
(1298),
(1296),
(1294),
(1292),
(1291),
(1289),
(1287),
(1286),
(1284),
(1282),
(1280),
(1279),
(1277),
(1275),
(1274),
(1272),
(1270),
(1269),
(1267),
(1265),
(1264),
(1262),
(1260),
(1259),
(1257),
(1256),
(1254),
(1252),
(1251),
(1249),
(1247),
(1246),
(1244),
(1243),
(1241),
(1239),
(1238),
(1236),
(1235),
(1233),
(1231),
(1230),
(1228),
(1227),
(1225),
(1224),
(1222),
(1221),
(1219),
(1218),
(1216),
(1214),
(1213),
(1211),
(1210),
(1208),
(1207),
(1205),
(1204),
(1202),
(1201),
(1199),
(1198),
(1196),
(1195),
(1193),
(1192),
(1190),
(1189),
(1187),
(1186),
(1185),
(1183),
(1182),
(1180),
(1179),
(1177),
(1176),
(1174),
(1173),
(1172),
(1170),
(1169),
(1167),
(1166),
(1164),
(1163),
(1162),
(1160),
(1159),
(1157),
(1156),
(1155),
(1153),
(1152),
(1151),
(1149),
(1148),
(1146),
(1145),
(1144),
(1142),
(1141),
(1140),
(1138),
(1137),
(1136),
(1134),
(1133),
(1132),
(1130),
(1129),
(1128),
(1126),
(1125),
(1124),
(1122),
(1121),
(1120),
(1118),
(1117),
(1116),
(1114),
(1113),
(1112),
(1111),
(1109),
(1108),
(1107),
(1105),
(1104),
(1103),
(1102),
(1100),
(1099),
(1098),
(1097),
(1095),
(1094),
(1093),
(1092),
(1090),
(1089),
(1088),
(1087),
(1085),
(1084),
(1083),
(1082),
(1080),
(1079),
(1078),
(1077),
(1076),
(1074),
(1073),
(1072),
(1071),
(1070),
(1068),
(1067),
(1066),
(1065),
(1064),
(1062),
(1061),
(1060),
(1059),
(1058),
(1057),
(1055),
(1054),
(1053),
(1052),
(1051),
(1050),
(1048),
(1047),
(1046),
(1045),
(1044),
(1043),
(1042),
(1040),
(1039),
(1038),
(1037),
(1036),
(1035),
(1034),
(1033),
(1031),
(1030),
(1029),
(1028),
(1027),
(1026),
(1025),
(1024),
(1023),
(1022),
(1020),
(1019),
(1018),
(1017),
(1016),
(1015),
(1014),
(1013),
(1012),
(1011),
(1010),
(1009),
(1007),
(1006),
(1005),
(1004),
(1003),
(1002),
(1001),
(1000),
(999),
(998),
(997),
(996),
(995),
(994),
(993),
(992),
(991),
(990),
(989),
(988),
(987),
(986),
(985),
(984),
(982),
(981),
(980),
(979),
(978),
(977),
(976),
(975),
(974),
(973),
(972),
(971),
(970),
(969),
(968),
(967),
(967),
(966),
(965),
(964),
(963),
(962),
(961),
(960),
(959),
(958),
(957),
(956),
(955),
(954),
(953),
(952),
(951),
(950),
(949),
(948),
(947),
(946),
(945),
(944),
(943),
(942),
(942),
(941),
(940),
(939),
(938),
(937),
(936),
(935),
(934),
(933),
(932),
(931),
(930),
(930),
(929),
(928),
(927),
(926),
(925),
(924),
(923),
(922),
(921),
(921),
(920),
(919),
(918),
(917),
(916),
(915),
(914),
(913),
(913),
(912),
(911),
(910),
(909),
(908),
(907),
(906),
(906),
(905),
(904),
(903),
(902),
(901),
(900),
(899),
(899),
(898),
(897),
(896),
(895),
(894),
(894),
(893),
(892),
(891),
(890),
(889),
(888),
(888),
(887),
(886),
(885),
(884),
(884),
(883),
(882),
(881),
(880),
(879),
(879),
(878),
(877),
(876),
(875),
(874),
(874),
(873),
(872),
(871),
(870),
(870),
(869),
(868),
(867),
(866),
(866),
(865),
(864),
(863),
(862),
(862),
(861),
(860),
(859),
(859),
(858),
(857),
(856),
(855),
(855),
(854),
(853),
(852),
(852),
(851),
(850),
(849),
(849),
(848),
(847),
(846),
(845),
(845),
(844),
(843),
(842),
(842),
(841),
(840),
(839),
(839),
(838),
(837),
(836),
(836),
(835),
(834),
(833),
(833),
(832),
(831),
(831),
(830),
(829),
(828),
(828),
(827),
(826),
(825),
(825),
(824),
(823),
(823),
(822),
(821),
(820),
(820),
(819),
(818),
(818),
(817),
(816),
(815),
(815),
(814),
(813),
(813),
(812),
(811),
(810),
(810),
(809),
(808),
(808),
(807),
(806),
(806),
(805),
(804),
(804),
(803),
(802),
(801),
(801),
(800),
(799),
(799),
(798),
(797),
(797),
(796),
(795),
(795),
(794),
(793),
(793),
(792),
(791),
(791),
(790),
(789),
(789),
(788),
(787),
(787),
(786),
(785),
(785),
(784),
(783),
(783),
(782),
(781),
(781),
(780),
(779),
(779),
(778),
(778),
(777),
(776),
(776),
(775),
(774),
(774),
(773),
(772),
(772),
(771),
(770),
(770),
(769),
(769),
(768),
(767),
(767),
(766),
(765),
(765),
(764),
(764),
(763),
(762),
(762),
(761),
(760),
(760),
(759),
(759),
(758),
(757),
(757),
(756),
(756),
(755),
(754),
(754),
(753),
(752),
(752),
(751),
(751),
(750),
(749),
(749),
(748),
(748),
(747),
(746),
(746),
(745),
(745),
(744),
(743),
(743),
(742),
(742),
(741),
(741),
(740),
(739),
(739),
(738),
(738),
(737),
(736),
(736),
(735),
(735),
(734),
(734),
(733),
(732),
(732),
(731),
(731),
(730),
(730),
(729),
(728),
(728),
(727),
(727),
(726),
(726),
(725),
(724),
(724),
(723),
(723),
(722),
(722),
(721),
(720),
(720),
(719),
(719),
(718),
(718),
(717),
(717),
(716),
(716),
(715),
(714),
(714),
(713),
(713),
(712),
(712),
(711),
(711),
(710),
(709),
(709),
(708),
(708),
(707),
(707),
(706),
(706),
(705),
(705),
(704),
(704),
(703),
(703),
(702),
(701),
(701),
(700),
(700),
(699),
(699),
(698),
(698),
(697),
(697),
(696),
(696),
(695),
(695),
(694),
(694),
(693),
(693),
(692),
(692),
(691),
(691),
(690),
(689),
(689),
(688),
(688),
(687),
(687),
(686),
(686),
(685),
(685),
(684),
(684),
(683),
(683),
(682),
(682),
(681),
(681),
(680),
(680),
(679),
(679),
(678),
(678),
(677),
(677),
(676),
(676),
(675),
(675),
(674),
(674),
(673),
(673),
(672),
(672),
(672),
(671),
(671),
(670),
(670),
(669),
(669),
(668),
(668),
(667),
(667),
(666),
(666),
(665),
(665),
(664),
(664),
(663),
(663),
(662),
(662),
(661),
(661),
(661),
(660),
(660),
(659),
(659),
(658),
(658),
(657),
(657),
(656),
(656),
(655),
(655),
(654),
(654),
(654),
(653),
(653),
(652),
(652),
(651),
(651),
(650),
(650),
(649),
(649),
(648),
(648),
(648),
(647),
(647),
(646),
(646),
(645),
(645),
(644),
(644),
(644),
(643),
(643),
(642),
(642),
(641),
(641),
(640),
(640),
(639),
(639),
(639),
(638),
(638),
(637),
(637),
(636),
(636),
(636),
(635),
(635),
(634),
(634),
(633),
(633),
(632),
(632),
(632),
(631),
(631),
(630),
(630),
(629),
(629),
(629),
(628),
(628),
(627),
(627),
(626),
(626),
(626),
(625),
(625),
(624),
(624),
(624),
(623),
(623),
(622),
(622),
(621),
(621),
(621),
(620),
(620),
(619),
(619),
(618),
(618),
(618),
(617),
(617),
(616),
(616),
(616),
(615),
(615),
(614),
(614),
(614),
(613),
(613),
(612),
(612),
(612),
(611),
(611),
(610),
(610),
(609),
(609),
(609),
(608),
(608),
(607),
(607),
(607),
(606),
(606),
(605),
(605),
(605),
(604),
(604),
(603),
(603),
(603),
(602),
(602),
(602),
(601),
(601),
(600),
(600),
(600),
(599),
(599),
(598),
(598),
(598),
(597),
(597),
(596),
(596),
(596),
(595),
(595),
(595),
(594),
(594),
(593),
(593),
(593),
(592),
(592),
(591),
(591),
(591),
(590),
(590),
(590),
(589),
(589),
(588),
(588),
(588),
(587),
(587),
(587),
(586),
(586),
(585),
(585),
(585),
(584),
(584),
(584),
(583),
(583),
(582),
(582),
(582),
(581),
(581),
(581),
(580),
(580),
(580),
(579),
(579),
(578),
(578),
(578),
(577),
(577),
(577),
(576),
(576),
(576),
(575),
(575),
(574),
(574),
(574),
(573),
(573),
(573),
(572),
(572),
(572),
(571),
(571),
(571),
(570),
(570),
(569),
(569),
(569),
(568),
(568),
(568),
(567),
(567),
(567),
(566),
(566),
(566),
(565),
(565),
(565),
(564),
(564),
(563),
(563),
(563),
(562),
(562),
(562),
(561),
(561),
(561),
(560),
(560),
(560),
(559),
(559),
(559),
(558),
(558),
(558),
(557),
(557),
(557),
(556),
(556),
(556),
(555),
(555),
(555),
(554),
(554),
(554),
(553),
(553),
(553),
(552),
(552),
(552),
(551),
(551),
(551),
(550),
(550),
(550),
(549),
(549),
(549),
(548),
(548),
(548),
(547),
(547),
(547),
(546),
(546),
(546),
(545),
(545),
(545),
(544),
(544),
(544),
(543),
(543),
(543),
(542),
(542),
(542),
(541),
(541),
(541),
(541),
(540),
(540),
(540),
(539),
(539),
(539),
(538),
(538),
(538),
(537),
(537),
(537),
(536),
(536),
(536),
(535),
(535),
(535),
(535),
(534),
(534),
(534),
(533),
(533),
(533),
(532),
(532),
(532),
(531),
(531),
(531),
(530),
(530),
(530),
(530),
(529),
(529),
(529),
(528),
(528),
(528),
(527),
(527),
(527),
(526),
(526),
(526),
(526),
(525),
(525),
(525),
(524),
(524),
(524),
(523),
(523),
(523),
(523),
(522),
(522),
(522),
(521),
(521),
(521),
(520),
(520),
(520),
(520),
(519),
(519),
(519),
(518),
(518),
(518),
(518),
(517),
(517),
(517),
(516),
(516),
(516),
(515),
(515),
(515),
(515),
(514),
(514),
(514),
(513),
(513),
(513),
(513),
(512),
(512),
(512),
(511),
(511),
(511),
(511),
(510),
(510),
(510),
(509),
(509),
(509),
(509),
(508),
(508),
(508),
(507),
(507),
(507),
(507),
(506),
(506),
(506),
(505),
(505),
(505),
(505),
(504),
(504),
(504),
(503),
(503),
(503),
(503),
(502),
(502),
(502),
(502),
(501),
(501),
(501),
(500),
(500),
(500),
(500),
(499),
(499),
(499),
(499),
(498),
(498),
(498),
(497),
(497),
(497),
(497),
(496),
(496),
(496),
(496),
(495),
(495),
(495),
(494),
(494),
(494),
(494),
(493),
(493),
(493),
(493),
(492),
(492),
(492),
(491),
(491),
(491),
(491),
(490),
(490),
(490),
(490),
(489),
(489),
(489),
(489),
(488),
(488),
(488),
(488),
(487),
(487),
(487),
(486),
(486),
(486),
(486),
(485),
(485),
(485),
(485),
(484),
(484),
(484),
(484),
(483),
(483),
(483),
(483),
(482),
(482),
(482),
(482),
(481),
(481),
(481),
(481),
(480),
(480),
(480),
(480),
(479),
(479),
(479),
(479),
(478),
(478),
(478),
(478),
(477),
(477),
(477),
(477),
(476),
(476),
(476),
(476),
(475),
(475),
(475),
(475),
(474),
(474),
(474),
(474),
(473),
(473),
(473),
(473),
(472),
(472),
(472),
(472),
(471),
(471),
(471),
(471),
(470),
(470),
(470),
(470),
(469),
(469),
(469),
(469),
(468),
(468),
(468),
(468),
(467),
(467),
(467),
(467),
(466),
(466),
(466),
(466),
(465),
(465),
(465),
(465),
(465),
(464),
(464),
(464),
(464),
(463),
(463),
(463),
(463),
(462),
(462),
(462),
(462),
(461),
(461),
(461),
(461),
(461),
(460),
(460),
(460),
(460),
(459),
(459),
(459),
(459),
(458),
(458),
(458),
(458),
(457),
(457),
(457),
(457),
(457),
(456),
(456),
(456),
(456),
(455),
(455),
(455),
(455),
(454),
(454),
(454),
(454),
(454),
(453),
(453),
(453),
(453),
(452),
(452),
(452),
(452),
(452),
(451),
(451),
(451),
(451),
(450),
(450),
(450),
(450),
(450),
(449),
(449),
(449),
(449),
(448),
(448),
(448),
(448),
(448),
(447),
(447),
(447),
(447),
(446),
(446),
(446),
(446),
(446),
(445),
(445),
(445),
(445),
(444),
(444),
(444),
(444),
(444),
(443),
(443),
(443),
(443),
(442),
(442),
(442),
(442),
(442),
(441),
(441),
(441),
(441),
(441),
(440),
(440),
(440),
(440),
(439),
(439),
(439),
(439),
(439),
(438),
(438),
(438),
(438),
(438),
(437),
(437),
(437),
(437),
(436),
(436),
(436),
(436),
(436),
(435),
(435),
(435),
(435),
(435),
(434),
(434),
(434),
(434),
(434),
(433),
(433),
(433),
(433),
(432),
(432),
(432),
(432),
(432),
(431),
(431),
(431),
(431),
(431),
(430),
(430),
(430),
(430),
(430),
(429),
(429),
(429),
(429),
(429),
(428),
(428),
(428),
(428),
(428),
(427),
(427),
(427),
(427),
(427),
(426),
(426),
(426),
(426),
(426),
(425),
(425),
(425),
(425),
(425),
(424),
(424),
(424),
(424),
(424),
(423),
(423),
(423),
(423),
(423),
(422),
(422),
(422),
(422),
(422),
(421),
(421),
(421),
(421),
(421),
(420),
(420),
(420),
(420),
(420),
(419),
(419),
(419),
(419),
(419),
(418),
(418),
(418),
(418),
(418),
(417),
(417),
(417),
(417),
(417),
(416),
(416),
(416),
(416),
(416),
(415),
(415),
(415),
(415),
(415),
(415),
(414),
(414),
(414),
(414),
(414),
(413),
(413),
(413),
(413),
(413),
(412),
(412),
(412),
(412),
(412),
(411),
(411),
(411),
(411),
(411),
(411),
(410),
(410),
(410),
(410),
(410),
(409),
(409),
(409),
(409),
(409),
(408),
(408),
(408),
(408),
(408),
(408),
(407),
(407),
(407),
(407),
(407),
(406),
(406),
(406),
(406),
(406),
(406),
(405),
(405),
(405),
(405),
(405),
(404),
(404),
(404),
(404),
(404),
(404),
(403),
(403),
(403),
(403),
(403),
(402),
(402),
(402),
(402),
(402),
(402),
(401),
(401),
(401),
(401),
(401),
(400),
(400),
(400),
(400),
(400),
(400),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0)

);


begin
		dist <= std_logic_vector(to_unsigned(table(to_integer(unsigned(volt))),dist'length));
		
end lookupTable;
	