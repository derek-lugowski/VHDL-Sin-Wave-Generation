library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity LUT_skip is 
	port(
		index		: in	std_logic_vector(11 downto 0);
		skip		: out	std_logic_vector(8 downto 0)
		);
end LUT_skip;

architecture lookupTable of LUT_skip is


type rom is array (0 to 4095) of integer;

constant table: rom:=(

(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(460),
(460),
(460),
(460),
(460),
(460),
(460),
(460),
(460),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468)


);


begin
		skip <= std_logic_vector(to_unsigned(table(to_integer(unsigned(index))),skip'length));
		
end lookupTable;
	