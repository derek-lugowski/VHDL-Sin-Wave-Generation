LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY sinval IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index          :  IN    STD_LOGIC_VECTOR(14 DOWNTO 0);-- change                           
      sin            :  OUT   STD_LOGIC_VECTOR(4 DOWNTO 0)); -- change 
END sinval;

ARCHITECTURE behavior OF sinval IS

-- multiplied sin value by 1023
-- skip by 468 for 650kHz

type array_1d is array (0 to 18000) of integer;
constant sin_LUT : array_1d := (
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(15),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(14),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(13),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(12),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(11),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(10),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(9),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(8),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(7),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(6),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(5),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(4),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(3),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(2),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(1),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0)


);


begin
    	
   sin <= std_logic_vector(to_unsigned(sin_LUT(to_integer(unsigned(index))),sin'length));

end behavior;